library verilog;
use verilog.vl_types.all;
entity mux_4to1_8b_test is
end mux_4to1_8b_test;
