library verilog;
use verilog.vl_types.all;
entity arithmeticMUX_test is
end arithmeticMUX_test;
