library verilog;
use verilog.vl_types.all;
entity fa_testbench is
end fa_testbench;
