library verilog;
use verilog.vl_types.all;
entity mux_4to1_1b_test is
end mux_4to1_1b_test;
