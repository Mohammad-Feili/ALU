library verilog;
use verilog.vl_types.all;
entity arithmeticU_test is
end arithmeticU_test;
