library verilog;
use verilog.vl_types.all;
entity LogicU_testbench is
end LogicU_testbench;
