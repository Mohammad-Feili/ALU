library verilog;
use verilog.vl_types.all;
entity arithmeticFA_test is
end arithmeticFA_test;
